module program_counter(
//inputs are target address of next instruction
//output is the instruction read from instruction mem
);

endmodule