module PCSrc (
//inputs include indicators that whether its a branch/jump/ret instruction
);

endmodule