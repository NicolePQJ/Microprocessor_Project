module dataMem(

);

endmodule