module REG(
//asynchronous write and synchronous read
);

endmodule