module insturction_mem(
//RISC-V instructions
);

endmodule